`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    12:07:22 03/02/2023 
// Design Name: 
// Module Name:    Gestor_de_perifricos 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module Gestor_de_perifricos(
    input ESCR_P,
    input [7:0] Operando1,
    input [7:0] PIN,
    output [7:0] Dados_IN,
    output [7:0] POUT
    );


endmodule
